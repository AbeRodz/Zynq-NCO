--------------------
-- SineLUT
-- Autor: Abraham R.
--------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity SineLUT is
  port (
    c_i    : in std_logic; -- Clock signal
    en_i   : in std_logic; -- Enable signal
    addr_i : in std_logic_vector(9 downto 0); -- Memory addres
    --
    wave_o : out std_logic_vector(15 downto 0) -- Output data
  );
end SineLUT;

architecture SineLUT_arq of SineLUT is

  type ROM is array (1023 downto 0) of integer range 0 to 65535; -- 10x16bit ROM

  signal t_ROM : ROM := (
  32767, 32968, 33169, 33370, 33571, 33772, 33973, 34174, 34375, 34576, 34776, 34977, 35177, 35378, 35578, 35779, 35979, 36179, 36379, 36578, 36778, 36977, 37177, 37376, 37575,
  37774, 37972, 38171, 38369, 38567, 38765, 38962, 39160, 39357, 39553, 39750, 39946, 40142, 40338, 40534, 40729, 40924, 41118, 41312, 41506, 41700, 41893, 42086, 42279, 42471,
  42663, 42854, 43045, 43236, 43426, 43616, 43806, 43995, 44184, 44372, 44560, 44747, 44934, 45120, 45306, 45492, 45677, 45861, 46046, 46229, 46412, 46595, 46777, 46958, 47139,
  47320, 47499, 47679, 47857, 48036, 48213, 48390, 48567, 48743, 48918, 49092, 49266, 49440, 49613, 49785, 49956, 50127, 50297, 50467, 50636, 50804, 50971, 51138, 51304, 51470,
  51635, 51799, 51962, 52124, 52286, 52447, 52608, 52767, 52926, 53084, 53242, 53398, 53554, 53709, 53863, 54017, 54170, 54321, 54472, 54623, 54772, 54921, 55068, 55215, 55361,
  55506, 55651, 55794, 55937, 56078, 56219, 56359, 56498, 56637, 56774, 56910, 57046, 57180, 57314, 57447, 57578, 57709, 57839, 57968, 58096, 58223, 58349, 58475, 58599, 58722,
  58844, 58965, 59086, 59205, 59323, 59441, 59557, 59672, 59786, 59900, 60012, 60123, 60233, 60342, 60450, 60557, 60663, 60768, 60872, 60975, 61077, 61178, 61277, 61376, 61473,
  61570, 61665, 61759, 61852, 61944, 62035, 62125, 62214, 62301, 62388, 62473, 62558, 62641, 62723, 62804, 62884, 62962, 63040, 63116, 63191, 63265, 63338, 63410, 63481, 63550,
  63619, 63686, 63752, 63817, 63880, 63943, 64004, 64064, 64123, 64181, 64237, 64293, 64347, 64400, 64452, 64503, 64552, 64600, 64647, 64693, 64738, 64781, 64824, 64865, 64904,
  64943, 64980, 65017, 65052, 65085, 65118, 65149, 65179, 65208, 65236, 65262, 65288, 65312, 65334, 65356, 65376, 65395, 65413, 65430, 65445, 65459, 65472, 65484, 65495, 65504,
  65512, 65519, 65524, 65528, 65532, 65533, 65534, 65533, 65532, 65528, 65524, 65519, 65512, 65504, 65495, 65484, 65472, 65459, 65445, 65430, 65413, 65395, 65376, 65356, 65334,
  65312, 65288, 65262, 65236, 65208, 65179, 65149, 65118, 65085, 65052, 65017, 64980, 64943, 64904, 64865, 64824, 64781, 64738, 64693, 64647, 64600, 64552, 64503, 64452, 64400,
  64347, 64293, 64237, 64181, 64123, 64064, 64004, 63943, 63880, 63817, 63752, 63686, 63619, 63550, 63481, 63410, 63338, 63265, 63191, 63116, 63040, 62962, 62884, 62804, 62723,
  62641, 62558, 62473, 62388, 62301, 62214, 62125, 62035, 61944, 61852, 61759, 61665, 61570, 61473, 61376, 61277, 61178, 61077, 60975, 60872, 60768, 60663, 60557, 60450, 60342,
  60233, 60123, 60012, 59900, 59786, 59672, 59557, 59441, 59323, 59205, 59086, 58965, 58844, 58722, 58599, 58475, 58349, 58223, 58096, 57968, 57839, 57709, 57578, 57447, 57314,
  57180, 57046, 56910, 56774, 56637, 56498, 56359, 56219, 56078, 55937, 55794, 55651, 55506, 55361, 55215, 55068, 54921, 54772, 54623, 54472, 54321, 54170, 54017, 53863, 53709,
  53554, 53398, 53242, 53084, 52926, 52767, 52608, 52447, 52286, 52124, 51962, 51799, 51635, 51470, 51304, 51138, 50971, 50804, 50636, 50467, 50297, 50127, 49956, 49785, 49613,
  49440, 49266, 49092, 48918, 48743, 48567, 48390, 48213, 48036, 47857, 47679, 47499, 47320, 47139, 46958, 46777, 46595, 46412, 46229, 46046, 45861, 45677, 45492, 45306, 45120,
  44934, 44747, 44560, 44372, 44184, 43995, 43806, 43616, 43426, 43236, 43045, 42854, 42663, 42471, 42279, 42086, 41893, 41700, 41506, 41312, 41118, 40924, 40729, 40534, 40338,
  40142, 39946, 39750, 39553, 39357, 39160, 38962, 38765, 38567, 38369, 38171, 37972, 37774, 37575, 37376, 37177, 36977, 36778, 36578, 36379, 36179, 35979, 35779, 35578, 35378,
  35177, 34977, 34776, 34576, 34375, 34174, 33973, 33772, 33571, 33370, 33169, 32968, 32767, 32566, 32365, 32164, 31963, 31762, 31561, 31360, 31159, 30958, 30758, 30557, 30357,
  30156, 29956, 29755, 29555, 29355, 29155, 28956, 28756, 28557, 28357, 28158, 27959, 27760, 27562, 27363, 27165, 26967, 26769, 26572, 26374, 26177, 25981, 25784, 25588, 25392,
  25196, 25000, 24805, 24610, 24416, 24222, 24028, 23834, 23641, 23448, 23255, 23063, 22871, 22680, 22489, 22298, 22108, 21918, 21728, 21539, 21350, 21162, 20974, 20787, 20600,
  20414, 20228, 20042, 19857, 19673, 19488, 19305, 19122, 18939, 18757, 18576, 18395, 18214, 18035, 17855, 17677, 17498, 17321, 17144, 16967, 16791, 16616, 16442, 16268, 16094,
  15921, 15749, 15578, 15407, 15237, 15067, 14898, 14730, 14563, 14396, 14230, 14064, 13899, 13735, 13572, 13410, 13248, 13087, 12926, 12767, 12608, 12450, 12292, 12136, 11980,
  11825, 11671, 11517, 11364, 11213, 11062, 10911, 10762, 10613, 10466, 10319, 10173, 10028, 9883, 9740, 9597, 9456, 9315, 9175, 9036, 8897, 8760, 8624, 8488, 8354,
  8220, 8087, 7956, 7825, 7695, 7566, 7438, 7311, 7185, 7059, 6935, 6812, 6690, 6569, 6448, 6329, 6211, 6093, 5977, 5862, 5748, 5634, 5522, 5411, 5301,
  5192, 5084, 4977, 4871, 4766, 4662, 4559, 4457, 4356, 4257, 4158, 4061, 3964, 3869, 3775, 3682, 3590, 3499, 3409, 3320, 3233, 3146, 3061, 2976, 2893,
  2811, 2730, 2650, 2572, 2494, 2418, 2343, 2269, 2196, 2124, 2053, 1984, 1915, 1848, 1782, 1717, 1654, 1591, 1530, 1470, 1411, 1353, 1297, 1241, 1187,
  1134, 1082, 1031, 982, 934, 887, 841, 796, 753, 710, 669, 630, 591, 554, 517, 482, 449, 416, 385, 355, 326, 298, 272, 246, 222,
  200, 178, 158, 139, 121, 104, 89, 75, 62, 50, 39, 30, 22, 15, 10, 6, 2, 1, 0, 1, 2, 6, 10, 15, 22,
  30, 39, 50, 62, 75, 89, 104, 121, 139, 158, 178, 200, 222, 246, 272, 298, 326, 355, 385, 416, 449, 482, 517, 554, 591,
  630, 669, 710, 753, 796, 841, 887, 934, 982, 1031, 1082, 1134, 1187, 1241, 1297, 1353, 1411, 1470, 1530, 1591, 1654, 1717, 1782, 1848, 1915,
  1984, 2053, 2124, 2196, 2269, 2343, 2418, 2494, 2572, 2650, 2730, 2811, 2893, 2976, 3061, 3146, 3233, 3320, 3409, 3499, 3590, 3682, 3775, 3869, 3964,
  4061, 4158, 4257, 4356, 4457, 4559, 4662, 4766, 4871, 4977, 5084, 5192, 5301, 5411, 5522, 5634, 5748, 5862, 5977, 6093, 6211, 6329, 6448, 6569, 6690,
  6812, 6935, 7059, 7185, 7311, 7438, 7566, 7695, 7825, 7956, 8087, 8220, 8354, 8488, 8624, 8760, 8897, 9036, 9175, 9315, 9456, 9597, 9740, 9883, 10028,
  10173, 10319, 10466, 10613, 10762, 10911, 11062, 11213, 11364, 11517, 11671, 11825, 11980, 12136, 12292, 12450, 12608, 12767, 12926, 13087, 13248, 13410, 13572, 13735, 13899,
  14064, 14230, 14396, 14563, 14730, 14898, 15067, 15237, 15407, 15578, 15749, 15921, 16094, 16268, 16442, 16616, 16791, 16967, 17144, 17321, 17498, 17677, 17855, 18035, 18214,
  18395, 18576, 18757, 18939, 19122, 19305, 19488, 19673, 19857, 20042, 20228, 20414, 20600, 20787, 20974, 21162, 21350, 21539, 21728, 21918, 22108, 22298, 22489, 22680, 22871,
  23063, 23255, 23448, 23641, 23834, 24028, 24222, 24416, 24610, 24805, 25000, 25196, 25392, 25588, 25784, 25981, 26177, 26374, 26572, 26769, 26967, 27165, 27363, 27562, 27760,
  27959, 28158, 28357, 28557, 28756, 28956, 29155, 29355, 29555, 29755, 29956, 30156, 30357, 30557, 30758, 30958, 31159, 31360, 31561, 31762, 31963, 32164, 32365, 32566

  );

begin

  SIN : process (c_i)
  begin
    if rising_edge(c_i) then
      if (en_i = '1') then
        wave_o <= std_logic_vector(to_Signed((t_ROM(to_Integer(Unsigned(addr_i))) - 32768), 16));
      end if;
    end if;
  end process SIN;

end;